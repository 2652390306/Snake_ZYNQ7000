module ctrl_game(
	input             lcd_pclk,     //ʱ��
    input             rst_n        //��λ���͵�ƽ��Ч
    );

endmodule
